`define NOP 2'b00 // No operation
`define MULTI 2'b11 // Mult imm and wait
`define ADDI 2'b01 // add immg